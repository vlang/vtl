module storage

import vtl.storage.vcl

// StorageDataType is a sum type that lists the possible types to be used to define storage
pub type StorageDataType = byte | f32 | f64 | i16 | i64 | i8 | int | u16 | u32 | u64

pub type Storage<T> = CpuStorage<T> | vcl.VclStorage<T>
