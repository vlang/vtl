module autograd


