module vtl
