module storage

fn test_cpu_with_default() {
	c := new_cpu_with_default(2, 0, int(sizeof(f64)), voidptr(0))
}
