module la

