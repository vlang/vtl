module vtl

pub const (
	version = '0.2'
)
