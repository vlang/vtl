module la
