module vnum

pub const (
	version = '0.1'
)
