module vtl


