module autograd
