module vtl

fn test_new() {
	t := new_tensor<f64>({
		shape: [3]
	})
}
