module la


